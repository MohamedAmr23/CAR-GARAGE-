library verilog;
use verilog.vl_types.all;
entity counter_g is
end counter_g;
