library verilog;
use verilog.vl_types.all;
entity clock_g is
end clock_g;
